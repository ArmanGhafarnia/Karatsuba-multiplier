LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;
USE ieee.std_logic_unsigned.ALL;
ENTITY loopback_Device IS
	PORT (
		nRST : IN STD_LOGIC;
		sys_clk : IN STD_LOGIC;
		nPause : IN STD_LOGIC;
		wren : OUT STD_LOGIC;
		tx_data : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		rx_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		rx_data_ready : IN STD_LOGIC;
		led_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		rx_data_accept : OUT STD_LOGIC;

		------------------------------------------------
		-- test vector signals should be configured 
		-- corresponding with the design
		-- Should be updated
		------------------------------------------------
		clk : OUT STD_LOGIC;
		rest : OUT STD_LOGIC;
		start : OUT STD_LOGIC;
		a : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
		b : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
		--
		p : IN STD_LOGIC_VECTOR(511 DOWNTO 0);
		done : IN STD_LOGIC
	);
END loopback_Device;

ARCHITECTURE behavioral OF loopback_Device IS
	----------------------------------------------------------------------
	-- Number of input and output bits: 
	-- Should be updated
	----------------------------------------------------------------------
	CONSTANT InputSize : INTEGER := 515; -- number of input bits
	CONSTANT OutputSize : INTEGER := 513; -- number of output bits
	----------------------------------------------------------------------
	CONSTANT CHAR0 : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00110000";
	CONSTANT CHAR1 : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00110001";
	TYPE reg_file IS ARRAY (0 TO 1030) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
	TYPE lp_state IS (wait_for_data, wait_one_cycle, send_output);

	SIGNAL state : lp_state;
	SIGNAL input_reg : reg_file;
	SIGNAL output_reg : reg_file;
	SIGNAL icntr, ocntr : INTEGER RANGE 0 TO 1030;
	SIGNAL dout : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL led_out_temp : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL led_out_cntr : STD_LOGIC_VECTOR(7 DOWNTO 0);
	FUNCTION c2s(x : STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
	BEGIN
		IF x = CHAR0 THEN
			RETURN '0';
		ELSE
			RETURN '1';
		END IF;
	END c2s;
	FUNCTION s2c(x : STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
	BEGIN
		IF x = '0' THEN
			RETURN CHAR0;
		ELSE
			RETURN CHAR1;
		END IF;
	END s2c;
BEGIN

	led_out <= led_out_cntr;

	seq : PROCESS (sys_clk, nRST)
	BEGIN
		IF nRST = '0' THEN
			tx_data <= (OTHERS => '0');
			wren <= '0';
			rx_data_accept <= '0';
			state <= wait_for_data;
			icntr <= 0;
			ocntr <= 0;
			led_out_temp <= (OTHERS => '0');
			led_out_cntr <= (OTHERS => '0');
		ELSIF sys_clk'EVENT AND sys_clk = '1' THEN
			IF nPause = '1' THEN
				wren <= '0';
				rx_data_accept <= '0';
				CASE state IS
					WHEN wait_for_data =>
						IF rx_data_ready = '1' THEN
							wren <= '1';
							rx_data_accept <= '1';
							IF icntr = InputSize THEN
								tx_data <= X"3D"; --=
								ocntr <= 0;
								state <= send_output;
							ELSE
								input_reg(icntr) <= rx_data;
								tx_data <= rx_data;
								icntr <= icntr + 1;
								state <= wait_one_cycle;
							END IF;
						END IF;
					WHEN wait_one_cycle =>
						rx_data_accept <= '0';
						wren <= '0';
						state <= wait_for_data;
					WHEN send_output =>
						wren <= '1';
						rx_data_accept <= '1';
						IF ocntr = OutputSize THEN
							tx_data <= X"23"; -- #
							state <= wait_one_cycle;
							icntr <= 0;
						ELSE
							tx_data <= output_reg(OutputSize - ocntr - 1);
							state <= send_output;
							ocntr <= ocntr + 1;
						END IF;
						led_out_cntr <= led_out_cntr + '1';
					WHEN OTHERS =>
						wren <= '0';
						rx_data_accept <= '0';
						tx_data <= (OTHERS => '0');
						tx_data <= rx_data;
						state <= wait_for_data;
				END CASE;
			END IF;
		END IF;
	END PROCESS seq;

	------------------------------------------
	-- Inteface with CUT: Should be updated
	-- Should be updated
	------------------------------------------

	-- convert input characters to bits
	clk <= c2s(input_reg(0));
	rest <= c2s(input_reg(1));
	start <= c2s(input_reg(2));
	a(255) <= c2s(input_reg(3));
	a(254) <= c2s(input_reg(4));
	a(253) <= c2s(input_reg(5));
	a(252) <= c2s(input_reg(6));
	a(251) <= c2s(input_reg(7));
	a(250) <= c2s(input_reg(8));
	a(249) <= c2s(input_reg(9));
	a(248) <= c2s(input_reg(10));
	a(247) <= c2s(input_reg(11));
	a(246) <= c2s(input_reg(12));
	a(245) <= c2s(input_reg(13));
	a(244) <= c2s(input_reg(14));
	a(243) <= c2s(input_reg(15));
	a(242) <= c2s(input_reg(16));
	a(241) <= c2s(input_reg(17));
	a(240) <= c2s(input_reg(18));
	a(239) <= c2s(input_reg(19));
	a(238) <= c2s(input_reg(20));
	a(237) <= c2s(input_reg(21));
	a(236) <= c2s(input_reg(22));
	a(235) <= c2s(input_reg(23));
	a(234) <= c2s(input_reg(24));
	a(233) <= c2s(input_reg(25));
	a(232) <= c2s(input_reg(26));
	a(231) <= c2s(input_reg(27));
	a(230) <= c2s(input_reg(28));
	a(229) <= c2s(input_reg(29));
	a(228) <= c2s(input_reg(30));
	a(227) <= c2s(input_reg(31));
	a(226) <= c2s(input_reg(32));
	a(225) <= c2s(input_reg(33));
	a(224) <= c2s(input_reg(34));
	a(223) <= c2s(input_reg(35));
	a(222) <= c2s(input_reg(36));
	a(221) <= c2s(input_reg(37));
	a(220) <= c2s(input_reg(38));
	a(219) <= c2s(input_reg(39));
	a(218) <= c2s(input_reg(40));
	a(217) <= c2s(input_reg(41));
	a(216) <= c2s(input_reg(42));
	a(215) <= c2s(input_reg(43));
	a(214) <= c2s(input_reg(44));
	a(213) <= c2s(input_reg(45));
	a(212) <= c2s(input_reg(46));
	a(211) <= c2s(input_reg(47));
	a(210) <= c2s(input_reg(48));
	a(209) <= c2s(input_reg(49));
	a(208) <= c2s(input_reg(50));
	a(207) <= c2s(input_reg(51));
	a(206) <= c2s(input_reg(52));
	a(205) <= c2s(input_reg(53));
	a(204) <= c2s(input_reg(54));
	a(203) <= c2s(input_reg(55));
	a(202) <= c2s(input_reg(56));
	a(201) <= c2s(input_reg(57));
	a(200) <= c2s(input_reg(58));
	a(199) <= c2s(input_reg(59));
	a(198) <= c2s(input_reg(60));
	a(197) <= c2s(input_reg(61));
	a(196) <= c2s(input_reg(62));
	a(195) <= c2s(input_reg(63));
	a(194) <= c2s(input_reg(64));
	a(193) <= c2s(input_reg(65));
	a(192) <= c2s(input_reg(66));
	a(191) <= c2s(input_reg(67));
	a(190) <= c2s(input_reg(68));
	a(189) <= c2s(input_reg(69));
	a(188) <= c2s(input_reg(70));
	a(187) <= c2s(input_reg(71));
	a(186) <= c2s(input_reg(72));
	a(185) <= c2s(input_reg(73));
	a(184) <= c2s(input_reg(74));
	a(183) <= c2s(input_reg(75));
	a(182) <= c2s(input_reg(76));
	a(181) <= c2s(input_reg(77));
	a(180) <= c2s(input_reg(78));
	a(179) <= c2s(input_reg(79));
	a(178) <= c2s(input_reg(80));
	a(177) <= c2s(input_reg(81));
	a(176) <= c2s(input_reg(82));
	a(175) <= c2s(input_reg(83));
	a(174) <= c2s(input_reg(84));
	a(173) <= c2s(input_reg(85));
	a(172) <= c2s(input_reg(86));
	a(171) <= c2s(input_reg(87));
	a(170) <= c2s(input_reg(88));
	a(169) <= c2s(input_reg(89));
	a(168) <= c2s(input_reg(90));
	a(167) <= c2s(input_reg(91));
	a(166) <= c2s(input_reg(92));
	a(165) <= c2s(input_reg(93));
	a(164) <= c2s(input_reg(94));
	a(163) <= c2s(input_reg(95));
	a(162) <= c2s(input_reg(96));
	a(161) <= c2s(input_reg(97));
	a(160) <= c2s(input_reg(98));
	a(159) <= c2s(input_reg(99));
	a(158) <= c2s(input_reg(100));
	a(157) <= c2s(input_reg(101));
	a(156) <= c2s(input_reg(102));
	a(155) <= c2s(input_reg(103));
	a(154) <= c2s(input_reg(104));
	a(153) <= c2s(input_reg(105));
	a(152) <= c2s(input_reg(106));
	a(151) <= c2s(input_reg(107));
	a(150) <= c2s(input_reg(108));
	a(149) <= c2s(input_reg(109));
	a(148) <= c2s(input_reg(110));
	a(147) <= c2s(input_reg(111));
	a(146) <= c2s(input_reg(112));
	a(145) <= c2s(input_reg(113));
	a(144) <= c2s(input_reg(114));
	a(143) <= c2s(input_reg(115));
	a(142) <= c2s(input_reg(116));
	a(141) <= c2s(input_reg(117));
	a(140) <= c2s(input_reg(118));
	a(139) <= c2s(input_reg(119));
	a(138) <= c2s(input_reg(120));
	a(137) <= c2s(input_reg(121));
	a(136) <= c2s(input_reg(122));
	a(135) <= c2s(input_reg(123));
	a(134) <= c2s(input_reg(124));
	a(133) <= c2s(input_reg(125));
	a(132) <= c2s(input_reg(126));
	a(131) <= c2s(input_reg(127));
	a(130) <= c2s(input_reg(128));
	a(129) <= c2s(input_reg(129));
	a(128) <= c2s(input_reg(130));
	a(127) <= c2s(input_reg(131));
	a(126) <= c2s(input_reg(132));
	a(125) <= c2s(input_reg(133));
	a(124) <= c2s(input_reg(134));
	a(123) <= c2s(input_reg(135));
	a(122) <= c2s(input_reg(136));
	a(121) <= c2s(input_reg(137));
	a(120) <= c2s(input_reg(138));
	a(119) <= c2s(input_reg(139));
	a(118) <= c2s(input_reg(140));
	a(117) <= c2s(input_reg(141));
	a(116) <= c2s(input_reg(142));
	a(115) <= c2s(input_reg(143));
	a(114) <= c2s(input_reg(144));
	a(113) <= c2s(input_reg(145));
	a(112) <= c2s(input_reg(146));
	a(111) <= c2s(input_reg(147));
	a(110) <= c2s(input_reg(148));
	a(109) <= c2s(input_reg(149));
	a(108) <= c2s(input_reg(150));
	a(107) <= c2s(input_reg(151));
	a(106) <= c2s(input_reg(152));
	a(105) <= c2s(input_reg(153));
	a(104) <= c2s(input_reg(154));
	a(103) <= c2s(input_reg(155));
	a(102) <= c2s(input_reg(156));
	a(101) <= c2s(input_reg(157));
	a(100) <= c2s(input_reg(158));
	a(99) <= c2s(input_reg(159));
	a(98) <= c2s(input_reg(160));
	a(97) <= c2s(input_reg(161));
	a(96) <= c2s(input_reg(162));
	a(95) <= c2s(input_reg(163));
	a(94) <= c2s(input_reg(164));
	a(93) <= c2s(input_reg(165));
	a(92) <= c2s(input_reg(166));
	a(91) <= c2s(input_reg(167));
	a(90) <= c2s(input_reg(168));
	a(89) <= c2s(input_reg(169));
	a(88) <= c2s(input_reg(170));
	a(87) <= c2s(input_reg(171));
	a(86) <= c2s(input_reg(172));
	a(85) <= c2s(input_reg(173));
	a(84) <= c2s(input_reg(174));
	a(83) <= c2s(input_reg(175));
	a(82) <= c2s(input_reg(176));
	a(81) <= c2s(input_reg(177));
	a(80) <= c2s(input_reg(178));
	a(79) <= c2s(input_reg(179));
	a(78) <= c2s(input_reg(180));
	a(77) <= c2s(input_reg(181));
	a(76) <= c2s(input_reg(182));
	a(75) <= c2s(input_reg(183));
	a(74) <= c2s(input_reg(184));
	a(73) <= c2s(input_reg(185));
	a(72) <= c2s(input_reg(186));
	a(71) <= c2s(input_reg(187));
	a(70) <= c2s(input_reg(188));
	a(69) <= c2s(input_reg(189));
	a(68) <= c2s(input_reg(190));
	a(67) <= c2s(input_reg(191));
	a(66) <= c2s(input_reg(192));
	a(65) <= c2s(input_reg(193));
	a(64) <= c2s(input_reg(194));
	a(63) <= c2s(input_reg(195));
	a(62) <= c2s(input_reg(196));
	a(61) <= c2s(input_reg(197));
	a(60) <= c2s(input_reg(198));
	a(59) <= c2s(input_reg(199));
	a(58) <= c2s(input_reg(200));
	a(57) <= c2s(input_reg(201));
	a(56) <= c2s(input_reg(202));
	a(55) <= c2s(input_reg(203));
	a(54) <= c2s(input_reg(204));
	a(53) <= c2s(input_reg(205));
	a(52) <= c2s(input_reg(206));
	a(51) <= c2s(input_reg(207));
	a(50) <= c2s(input_reg(208));
	a(49) <= c2s(input_reg(209));
	a(48) <= c2s(input_reg(210));
	a(47) <= c2s(input_reg(211));
	a(46) <= c2s(input_reg(212));
	a(45) <= c2s(input_reg(213));
	a(44) <= c2s(input_reg(214));
	a(43) <= c2s(input_reg(215));
	a(42) <= c2s(input_reg(216));
	a(41) <= c2s(input_reg(217));
	a(40) <= c2s(input_reg(218));
	a(39) <= c2s(input_reg(219));
	a(38) <= c2s(input_reg(220));
	a(37) <= c2s(input_reg(221));
	a(36) <= c2s(input_reg(222));
	a(35) <= c2s(input_reg(223));
	a(34) <= c2s(input_reg(224));
	a(33) <= c2s(input_reg(225));
	a(32) <= c2s(input_reg(226));
	a(31) <= c2s(input_reg(227));
	a(30) <= c2s(input_reg(228));
	a(29) <= c2s(input_reg(229));
	a(28) <= c2s(input_reg(230));
	a(27) <= c2s(input_reg(231));
	a(26) <= c2s(input_reg(232));
	a(25) <= c2s(input_reg(233));
	a(24) <= c2s(input_reg(234));
	a(23) <= c2s(input_reg(235));
	a(22) <= c2s(input_reg(236));
	a(21) <= c2s(input_reg(237));
	a(20) <= c2s(input_reg(238));
	a(19) <= c2s(input_reg(239));
	a(18) <= c2s(input_reg(240));
	a(17) <= c2s(input_reg(241));
	a(16) <= c2s(input_reg(242));
	a(15) <= c2s(input_reg(243));
	a(14) <= c2s(input_reg(244));
	a(13) <= c2s(input_reg(245));
	a(12) <= c2s(input_reg(246));
	a(11) <= c2s(input_reg(247));
	a(10) <= c2s(input_reg(248));
	a(9) <= c2s(input_reg(249));
	a(8) <= c2s(input_reg(250));
	a(7) <= c2s(input_reg(251));
	a(6) <= c2s(input_reg(252));
	a(5) <= c2s(input_reg(253));
	a(4) <= c2s(input_reg(254));
	a(3) <= c2s(input_reg(255));
	a(2) <= c2s(input_reg(256));
	a(1) <= c2s(input_reg(257));
	a(0) <= c2s(input_reg(258));
	b(255) <= c2s(input_reg(259));
	b(254) <= c2s(input_reg(260));
	b(253) <= c2s(input_reg(261));
	b(252) <= c2s(input_reg(262));
	b(251) <= c2s(input_reg(263));
	b(250) <= c2s(input_reg(264));
	b(249) <= c2s(input_reg(265));
	b(248) <= c2s(input_reg(266));
	b(247) <= c2s(input_reg(267));
	b(246) <= c2s(input_reg(268));
	b(245) <= c2s(input_reg(269));
	b(244) <= c2s(input_reg(270));
	b(243) <= c2s(input_reg(271));
	b(242) <= c2s(input_reg(272));
	b(241) <= c2s(input_reg(273));
	b(240) <= c2s(input_reg(274));
	b(239) <= c2s(input_reg(275));
	b(238) <= c2s(input_reg(276));
	b(237) <= c2s(input_reg(277));
	b(236) <= c2s(input_reg(278));
	b(235) <= c2s(input_reg(279));
	b(234) <= c2s(input_reg(280));
	b(233) <= c2s(input_reg(281));
	b(232) <= c2s(input_reg(282));
	b(231) <= c2s(input_reg(283));
	b(230) <= c2s(input_reg(284));
	b(229) <= c2s(input_reg(285));
	b(228) <= c2s(input_reg(286));
	b(227) <= c2s(input_reg(287));
	b(226) <= c2s(input_reg(288));
	b(225) <= c2s(input_reg(289));
	b(224) <= c2s(input_reg(290));
	b(223) <= c2s(input_reg(291));
	b(222) <= c2s(input_reg(292));
	b(221) <= c2s(input_reg(293));
	b(220) <= c2s(input_reg(294));
	b(219) <= c2s(input_reg(295));
	b(218) <= c2s(input_reg(296));
	b(217) <= c2s(input_reg(297));
	b(216) <= c2s(input_reg(298));
	b(215) <= c2s(input_reg(299));
	b(214) <= c2s(input_reg(300));
	b(213) <= c2s(input_reg(301));
	b(212) <= c2s(input_reg(302));
	b(211) <= c2s(input_reg(303));
	b(210) <= c2s(input_reg(304));
	b(209) <= c2s(input_reg(305));
	b(208) <= c2s(input_reg(306));
	b(207) <= c2s(input_reg(307));
	b(206) <= c2s(input_reg(308));
	b(205) <= c2s(input_reg(309));
	b(204) <= c2s(input_reg(310));
	b(203) <= c2s(input_reg(311));
	b(202) <= c2s(input_reg(312));
	b(201) <= c2s(input_reg(313));
	b(200) <= c2s(input_reg(314));
	b(199) <= c2s(input_reg(315));
	b(198) <= c2s(input_reg(316));
	b(197) <= c2s(input_reg(317));
	b(196) <= c2s(input_reg(318));
	b(195) <= c2s(input_reg(319));
	b(194) <= c2s(input_reg(320));
	b(193) <= c2s(input_reg(321));
	b(192) <= c2s(input_reg(322));
	b(191) <= c2s(input_reg(323));
	b(190) <= c2s(input_reg(324));
	b(189) <= c2s(input_reg(325));
	b(188) <= c2s(input_reg(326));
	b(187) <= c2s(input_reg(327));
	b(186) <= c2s(input_reg(328));
	b(185) <= c2s(input_reg(329));
	b(184) <= c2s(input_reg(330));
	b(183) <= c2s(input_reg(331));
	b(182) <= c2s(input_reg(332));
	b(181) <= c2s(input_reg(333));
	b(180) <= c2s(input_reg(334));
	b(179) <= c2s(input_reg(335));
	b(178) <= c2s(input_reg(336));
	b(177) <= c2s(input_reg(337));
	b(176) <= c2s(input_reg(338));
	b(175) <= c2s(input_reg(339));
	b(174) <= c2s(input_reg(340));
	b(173) <= c2s(input_reg(341));
	b(172) <= c2s(input_reg(342));
	b(171) <= c2s(input_reg(343));
	b(170) <= c2s(input_reg(344));
	b(169) <= c2s(input_reg(345));
	b(168) <= c2s(input_reg(346));
	b(167) <= c2s(input_reg(347));
	b(166) <= c2s(input_reg(348));
	b(165) <= c2s(input_reg(349));
	b(164) <= c2s(input_reg(350));
	b(163) <= c2s(input_reg(351));
	b(162) <= c2s(input_reg(352));
	b(161) <= c2s(input_reg(353));
	b(160) <= c2s(input_reg(354));
	b(159) <= c2s(input_reg(355));
	b(158) <= c2s(input_reg(356));
	b(157) <= c2s(input_reg(357));
	b(156) <= c2s(input_reg(358));
	b(155) <= c2s(input_reg(359));
	b(154) <= c2s(input_reg(360));
	b(153) <= c2s(input_reg(361));
	b(152) <= c2s(input_reg(362));
	b(151) <= c2s(input_reg(363));
	b(150) <= c2s(input_reg(364));
	b(149) <= c2s(input_reg(365));
	b(148) <= c2s(input_reg(366));
	b(147) <= c2s(input_reg(367));
	b(146) <= c2s(input_reg(368));
	b(145) <= c2s(input_reg(369));
	b(144) <= c2s(input_reg(370));
	b(143) <= c2s(input_reg(371));
	b(142) <= c2s(input_reg(372));
	b(141) <= c2s(input_reg(373));
	b(140) <= c2s(input_reg(374));
	b(139) <= c2s(input_reg(375));
	b(138) <= c2s(input_reg(376));
	b(137) <= c2s(input_reg(377));
	b(136) <= c2s(input_reg(378));
	b(135) <= c2s(input_reg(379));
	b(134) <= c2s(input_reg(380));
	b(133) <= c2s(input_reg(381));
	b(132) <= c2s(input_reg(382));
	b(131) <= c2s(input_reg(383));
	b(130) <= c2s(input_reg(384));
	b(129) <= c2s(input_reg(385));
	b(128) <= c2s(input_reg(386));
	b(127) <= c2s(input_reg(387));
	b(126) <= c2s(input_reg(388));
	b(125) <= c2s(input_reg(389));
	b(124) <= c2s(input_reg(390));
	b(123) <= c2s(input_reg(391));
	b(122) <= c2s(input_reg(392));
	b(121) <= c2s(input_reg(393));
	b(120) <= c2s(input_reg(394));
	b(119) <= c2s(input_reg(395));
	b(118) <= c2s(input_reg(396));
	b(117) <= c2s(input_reg(397));
	b(116) <= c2s(input_reg(398));
	b(115) <= c2s(input_reg(399));
	b(114) <= c2s(input_reg(400));
	b(113) <= c2s(input_reg(401));
	b(112) <= c2s(input_reg(402));
	b(111) <= c2s(input_reg(403));
	b(110) <= c2s(input_reg(404));
	b(109) <= c2s(input_reg(405));
	b(108) <= c2s(input_reg(406));
	b(107) <= c2s(input_reg(407));
	b(106) <= c2s(input_reg(408));
	b(105) <= c2s(input_reg(409));
	b(104) <= c2s(input_reg(410));
	b(103) <= c2s(input_reg(411));
	b(102) <= c2s(input_reg(412));
	b(101) <= c2s(input_reg(413));
	b(100) <= c2s(input_reg(414));
	b(99) <= c2s(input_reg(415));
	b(98) <= c2s(input_reg(416));
	b(97) <= c2s(input_reg(417));
	b(96) <= c2s(input_reg(418));
	b(95) <= c2s(input_reg(419));
	b(94) <= c2s(input_reg(420));
	b(93) <= c2s(input_reg(421));
	b(92) <= c2s(input_reg(422));
	b(91) <= c2s(input_reg(423));
	b(90) <= c2s(input_reg(424));
	b(89) <= c2s(input_reg(425));
	b(88) <= c2s(input_reg(426));
	b(87) <= c2s(input_reg(427));
	b(86) <= c2s(input_reg(428));
	b(85) <= c2s(input_reg(429));
	b(84) <= c2s(input_reg(430));
	b(83) <= c2s(input_reg(431));
	b(82) <= c2s(input_reg(432));
	b(81) <= c2s(input_reg(433));
	b(80) <= c2s(input_reg(434));
	b(79) <= c2s(input_reg(435));
	b(78) <= c2s(input_reg(436));
	b(77) <= c2s(input_reg(437));
	b(76) <= c2s(input_reg(438));
	b(75) <= c2s(input_reg(439));
	b(74) <= c2s(input_reg(440));
	b(73) <= c2s(input_reg(441));
	b(72) <= c2s(input_reg(442));
	b(71) <= c2s(input_reg(443));
	b(70) <= c2s(input_reg(444));
	b(69) <= c2s(input_reg(445));
	b(68) <= c2s(input_reg(446));
	b(67) <= c2s(input_reg(447));
	b(66) <= c2s(input_reg(448));
	b(65) <= c2s(input_reg(449));
	b(64) <= c2s(input_reg(450));
	b(63) <= c2s(input_reg(451));
	b(62) <= c2s(input_reg(452));
	b(61) <= c2s(input_reg(453));
	b(60) <= c2s(input_reg(454));
	b(59) <= c2s(input_reg(455));
	b(58) <= c2s(input_reg(456));
	b(57) <= c2s(input_reg(457));
	b(56) <= c2s(input_reg(458));
	b(55) <= c2s(input_reg(459));
	b(54) <= c2s(input_reg(460));
	b(53) <= c2s(input_reg(461));
	b(52) <= c2s(input_reg(462));
	b(51) <= c2s(input_reg(463));
	b(50) <= c2s(input_reg(464));
	b(49) <= c2s(input_reg(465));
	b(48) <= c2s(input_reg(466));
	b(47) <= c2s(input_reg(467));
	b(46) <= c2s(input_reg(468));
	b(45) <= c2s(input_reg(469));
	b(44) <= c2s(input_reg(470));
	b(43) <= c2s(input_reg(471));
	b(42) <= c2s(input_reg(472));
	b(41) <= c2s(input_reg(473));
	b(40) <= c2s(input_reg(474));
	b(39) <= c2s(input_reg(475));
	b(38) <= c2s(input_reg(476));
	b(37) <= c2s(input_reg(477));
	b(36) <= c2s(input_reg(478));
	b(35) <= c2s(input_reg(479));
	b(34) <= c2s(input_reg(480));
	b(33) <= c2s(input_reg(481));
	b(32) <= c2s(input_reg(482));
	b(31) <= c2s(input_reg(483));
	b(30) <= c2s(input_reg(484));
	b(29) <= c2s(input_reg(485));
	b(28) <= c2s(input_reg(486));
	b(27) <= c2s(input_reg(487));
	b(26) <= c2s(input_reg(488));
	b(25) <= c2s(input_reg(489));
	b(24) <= c2s(input_reg(490));
	b(23) <= c2s(input_reg(491));
	b(22) <= c2s(input_reg(492));
	b(21) <= c2s(input_reg(493));
	b(20) <= c2s(input_reg(494));
	b(19) <= c2s(input_reg(495));
	b(18) <= c2s(input_reg(496));
	b(17) <= c2s(input_reg(497));
	b(16) <= c2s(input_reg(498));
	b(15) <= c2s(input_reg(499));
	b(14) <= c2s(input_reg(500));
	b(13) <= c2s(input_reg(501));
	b(12) <= c2s(input_reg(502));
	b(11) <= c2s(input_reg(503));
	b(10) <= c2s(input_reg(504));
	b(9) <= c2s(input_reg(505));
	b(8) <= c2s(input_reg(506));
	b(7) <= c2s(input_reg(507));
	b(6) <= c2s(input_reg(508));
	b(5) <= c2s(input_reg(509));
	b(4) <= c2s(input_reg(510));
	b(3) <= c2s(input_reg(511));
	b(2) <= c2s(input_reg(512));
	b(1) <= c2s(input_reg(513));
	b(0) <= c2s(input_reg(514));
	
	-- convert output bits to character
	output_reg(512) <= s2c(p(511));
	output_reg(511) <= s2c(p(510));
	output_reg(510) <= s2c(p(509));
	output_reg(509) <= s2c(p(508));
	output_reg(508) <= s2c(p(507));
	output_reg(507) <= s2c(p(506));
	output_reg(506) <= s2c(p(505));
	output_reg(505) <= s2c(p(504));
	output_reg(504) <= s2c(p(503));
	output_reg(503) <= s2c(p(502));
	output_reg(502) <= s2c(p(501));
	output_reg(501) <= s2c(p(500));
	output_reg(500) <= s2c(p(499));
	output_reg(499) <= s2c(p(498));
	output_reg(498) <= s2c(p(497));
	output_reg(497) <= s2c(p(496));
	output_reg(496) <= s2c(p(495));
	output_reg(495) <= s2c(p(494));
	output_reg(494) <= s2c(p(493));
	output_reg(493) <= s2c(p(492));
	output_reg(492) <= s2c(p(491));
	output_reg(491) <= s2c(p(490));
	output_reg(490) <= s2c(p(489));
	output_reg(489) <= s2c(p(488));
	output_reg(488) <= s2c(p(487));
	output_reg(487) <= s2c(p(486));
	output_reg(486) <= s2c(p(485));
	output_reg(485) <= s2c(p(484));
	output_reg(484) <= s2c(p(483));
	output_reg(483) <= s2c(p(482));
	output_reg(482) <= s2c(p(481));
	output_reg(481) <= s2c(p(480));
	output_reg(480) <= s2c(p(479));
	output_reg(479) <= s2c(p(478));
	output_reg(478) <= s2c(p(477));
	output_reg(477) <= s2c(p(476));
	output_reg(476) <= s2c(p(475));
	output_reg(475) <= s2c(p(474));
	output_reg(474) <= s2c(p(473));
	output_reg(473) <= s2c(p(472));
	output_reg(472) <= s2c(p(471));
	output_reg(471) <= s2c(p(470));
	output_reg(470) <= s2c(p(469));
	output_reg(469) <= s2c(p(468));
	output_reg(468) <= s2c(p(467));
	output_reg(467) <= s2c(p(466));
	output_reg(466) <= s2c(p(465));
	output_reg(465) <= s2c(p(464));
	output_reg(464) <= s2c(p(463));
	output_reg(463) <= s2c(p(462));
	output_reg(462) <= s2c(p(461));
	output_reg(461) <= s2c(p(460));
	output_reg(460) <= s2c(p(459));
	output_reg(459) <= s2c(p(458));
	output_reg(458) <= s2c(p(457));
	output_reg(457) <= s2c(p(456));
	output_reg(456) <= s2c(p(455));
	output_reg(455) <= s2c(p(454));
	output_reg(454) <= s2c(p(453));
	output_reg(453) <= s2c(p(452));
	output_reg(452) <= s2c(p(451));
	output_reg(451) <= s2c(p(450));
	output_reg(450) <= s2c(p(449));
	output_reg(449) <= s2c(p(448));
	output_reg(448) <= s2c(p(447));
	output_reg(447) <= s2c(p(446));
	output_reg(446) <= s2c(p(445));
	output_reg(445) <= s2c(p(444));
	output_reg(444) <= s2c(p(443));
	output_reg(443) <= s2c(p(442));
	output_reg(442) <= s2c(p(441));
	output_reg(441) <= s2c(p(440));
	output_reg(440) <= s2c(p(439));
	output_reg(439) <= s2c(p(438));
	output_reg(438) <= s2c(p(437));
	output_reg(437) <= s2c(p(436));
	output_reg(436) <= s2c(p(435));
	output_reg(435) <= s2c(p(434));
	output_reg(434) <= s2c(p(433));
	output_reg(433) <= s2c(p(432));
	output_reg(432) <= s2c(p(431));
	output_reg(431) <= s2c(p(430));
	output_reg(430) <= s2c(p(429));
	output_reg(429) <= s2c(p(428));
	output_reg(428) <= s2c(p(427));
	output_reg(427) <= s2c(p(426));
	output_reg(426) <= s2c(p(425));
	output_reg(425) <= s2c(p(424));
	output_reg(424) <= s2c(p(423));
	output_reg(423) <= s2c(p(422));
	output_reg(422) <= s2c(p(421));
	output_reg(421) <= s2c(p(420));
	output_reg(420) <= s2c(p(419));
	output_reg(419) <= s2c(p(418));
	output_reg(418) <= s2c(p(417));
	output_reg(417) <= s2c(p(416));
	output_reg(416) <= s2c(p(415));
	output_reg(415) <= s2c(p(414));
	output_reg(414) <= s2c(p(413));
	output_reg(413) <= s2c(p(412));
	output_reg(412) <= s2c(p(411));
	output_reg(411) <= s2c(p(410));
	output_reg(410) <= s2c(p(409));
	output_reg(409) <= s2c(p(408));
	output_reg(408) <= s2c(p(407));
	output_reg(407) <= s2c(p(406));
	output_reg(406) <= s2c(p(405));
	output_reg(405) <= s2c(p(404));
	output_reg(404) <= s2c(p(403));
	output_reg(403) <= s2c(p(402));
	output_reg(402) <= s2c(p(401));
	output_reg(401) <= s2c(p(400));
	output_reg(400) <= s2c(p(399));
	output_reg(399) <= s2c(p(398));
	output_reg(398) <= s2c(p(397));
	output_reg(397) <= s2c(p(396));
	output_reg(396) <= s2c(p(395));
	output_reg(395) <= s2c(p(394));
	output_reg(394) <= s2c(p(393));
	output_reg(393) <= s2c(p(392));
	output_reg(392) <= s2c(p(391));
	output_reg(391) <= s2c(p(390));
	output_reg(390) <= s2c(p(389));
	output_reg(389) <= s2c(p(388));
	output_reg(388) <= s2c(p(387));
	output_reg(387) <= s2c(p(386));
	output_reg(386) <= s2c(p(385));
	output_reg(385) <= s2c(p(384));
	output_reg(384) <= s2c(p(383));
	output_reg(383) <= s2c(p(382));
	output_reg(382) <= s2c(p(381));
	output_reg(381) <= s2c(p(380));
	output_reg(380) <= s2c(p(379));
	output_reg(379) <= s2c(p(378));
	output_reg(378) <= s2c(p(377));
	output_reg(377) <= s2c(p(376));
	output_reg(376) <= s2c(p(375));
	output_reg(375) <= s2c(p(374));
	output_reg(374) <= s2c(p(373));
	output_reg(373) <= s2c(p(372));
	output_reg(372) <= s2c(p(371));
	output_reg(371) <= s2c(p(370));
	output_reg(370) <= s2c(p(369));
	output_reg(369) <= s2c(p(368));
	output_reg(368) <= s2c(p(367));
	output_reg(367) <= s2c(p(366));
	output_reg(366) <= s2c(p(365));
	output_reg(365) <= s2c(p(364));
	output_reg(364) <= s2c(p(363));
	output_reg(363) <= s2c(p(362));
	output_reg(362) <= s2c(p(361));
	output_reg(361) <= s2c(p(360));
	output_reg(360) <= s2c(p(359));
	output_reg(359) <= s2c(p(358));
	output_reg(358) <= s2c(p(357));
	output_reg(357) <= s2c(p(356));
	output_reg(356) <= s2c(p(355));
	output_reg(355) <= s2c(p(354));
	output_reg(354) <= s2c(p(353));
	output_reg(353) <= s2c(p(352));
	output_reg(352) <= s2c(p(351));
	output_reg(351) <= s2c(p(350));
	output_reg(350) <= s2c(p(349));
	output_reg(349) <= s2c(p(348));
	output_reg(348) <= s2c(p(347));
	output_reg(347) <= s2c(p(346));
	output_reg(346) <= s2c(p(345));
	output_reg(345) <= s2c(p(344));
	output_reg(344) <= s2c(p(343));
	output_reg(343) <= s2c(p(342));
	output_reg(342) <= s2c(p(341));
	output_reg(341) <= s2c(p(340));
	output_reg(340) <= s2c(p(339));
	output_reg(339) <= s2c(p(338));
	output_reg(338) <= s2c(p(337));
	output_reg(337) <= s2c(p(336));
	output_reg(336) <= s2c(p(335));
	output_reg(335) <= s2c(p(334));
	output_reg(334) <= s2c(p(333));
	output_reg(333) <= s2c(p(332));
	output_reg(332) <= s2c(p(331));
	output_reg(331) <= s2c(p(330));
	output_reg(330) <= s2c(p(329));
	output_reg(329) <= s2c(p(328));
	output_reg(328) <= s2c(p(327));
	output_reg(327) <= s2c(p(326));
	output_reg(326) <= s2c(p(325));
	output_reg(325) <= s2c(p(324));
	output_reg(324) <= s2c(p(323));
	output_reg(323) <= s2c(p(322));
	output_reg(322) <= s2c(p(321));
	output_reg(321) <= s2c(p(320));
	output_reg(320) <= s2c(p(319));
	output_reg(319) <= s2c(p(318));
	output_reg(318) <= s2c(p(317));
	output_reg(317) <= s2c(p(316));
	output_reg(316) <= s2c(p(315));
	output_reg(315) <= s2c(p(314));
	output_reg(314) <= s2c(p(313));
	output_reg(313) <= s2c(p(312));
	output_reg(312) <= s2c(p(311));
	output_reg(311) <= s2c(p(310));
	output_reg(310) <= s2c(p(309));
	output_reg(309) <= s2c(p(308));
	output_reg(308) <= s2c(p(307));
	output_reg(307) <= s2c(p(306));
	output_reg(306) <= s2c(p(305));
	output_reg(305) <= s2c(p(304));
	output_reg(304) <= s2c(p(303));
	output_reg(303) <= s2c(p(302));
	output_reg(302) <= s2c(p(301));
	output_reg(301) <= s2c(p(300));
	output_reg(300) <= s2c(p(299));
	output_reg(299) <= s2c(p(298));
	output_reg(298) <= s2c(p(297));
	output_reg(297) <= s2c(p(296));
	output_reg(296) <= s2c(p(295));
	output_reg(295) <= s2c(p(294));
	output_reg(294) <= s2c(p(293));
	output_reg(293) <= s2c(p(292));
	output_reg(292) <= s2c(p(291));
	output_reg(291) <= s2c(p(290));
	output_reg(290) <= s2c(p(289));
	output_reg(289) <= s2c(p(288));
	output_reg(288) <= s2c(p(287));
	output_reg(287) <= s2c(p(286));
	output_reg(286) <= s2c(p(285));
	output_reg(285) <= s2c(p(284));
	output_reg(284) <= s2c(p(283));
	output_reg(283) <= s2c(p(282));
	output_reg(282) <= s2c(p(281));
	output_reg(281) <= s2c(p(280));
	output_reg(280) <= s2c(p(279));
	output_reg(279) <= s2c(p(278));
	output_reg(278) <= s2c(p(277));
	output_reg(277) <= s2c(p(276));
	output_reg(276) <= s2c(p(275));
	output_reg(275) <= s2c(p(274));
	output_reg(274) <= s2c(p(273));
	output_reg(273) <= s2c(p(272));
	output_reg(272) <= s2c(p(271));
	output_reg(271) <= s2c(p(270));
	output_reg(270) <= s2c(p(269));
	output_reg(269) <= s2c(p(268));
	output_reg(268) <= s2c(p(267));
	output_reg(267) <= s2c(p(266));
	output_reg(266) <= s2c(p(265));
	output_reg(265) <= s2c(p(264));
	output_reg(264) <= s2c(p(263));
	output_reg(263) <= s2c(p(262));
	output_reg(262) <= s2c(p(261));
	output_reg(261) <= s2c(p(260));
	output_reg(260) <= s2c(p(259));
	output_reg(259) <= s2c(p(258));
	output_reg(258) <= s2c(p(257));
	output_reg(257) <= s2c(p(256));
	output_reg(256) <= s2c(p(255));
	output_reg(255) <= s2c(p(254));
	output_reg(254) <= s2c(p(253));
	output_reg(253) <= s2c(p(252));
	output_reg(252) <= s2c(p(251));
	output_reg(251) <= s2c(p(250));
	output_reg(250) <= s2c(p(249));
	output_reg(249) <= s2c(p(248));
	output_reg(248) <= s2c(p(247));
	output_reg(247) <= s2c(p(246));
	output_reg(246) <= s2c(p(245));
	output_reg(245) <= s2c(p(244));
	output_reg(244) <= s2c(p(243));
	output_reg(243) <= s2c(p(242));
	output_reg(242) <= s2c(p(241));
	output_reg(241) <= s2c(p(240));
	output_reg(240) <= s2c(p(239));
	output_reg(239) <= s2c(p(238));
	output_reg(238) <= s2c(p(237));
	output_reg(237) <= s2c(p(236));
	output_reg(236) <= s2c(p(235));
	output_reg(235) <= s2c(p(234));
	output_reg(234) <= s2c(p(233));
	output_reg(233) <= s2c(p(232));
	output_reg(232) <= s2c(p(231));
	output_reg(231) <= s2c(p(230));
	output_reg(230) <= s2c(p(229));
	output_reg(229) <= s2c(p(228));
	output_reg(228) <= s2c(p(227));
	output_reg(227) <= s2c(p(226));
	output_reg(226) <= s2c(p(225));
	output_reg(225) <= s2c(p(224));
	output_reg(224) <= s2c(p(223));
	output_reg(223) <= s2c(p(222));
	output_reg(222) <= s2c(p(221));
	output_reg(221) <= s2c(p(220));
	output_reg(220) <= s2c(p(219));
	output_reg(219) <= s2c(p(218));
	output_reg(218) <= s2c(p(217));
	output_reg(217) <= s2c(p(216));
	output_reg(216) <= s2c(p(215));
	output_reg(215) <= s2c(p(214));
	output_reg(214) <= s2c(p(213));
	output_reg(213) <= s2c(p(212));
	output_reg(212) <= s2c(p(211));
	output_reg(211) <= s2c(p(210));
	output_reg(210) <= s2c(p(209));
	output_reg(209) <= s2c(p(208));
	output_reg(208) <= s2c(p(207));
	output_reg(207) <= s2c(p(206));
	output_reg(206) <= s2c(p(205));
	output_reg(205) <= s2c(p(204));
	output_reg(204) <= s2c(p(203));
	output_reg(203) <= s2c(p(202));
	output_reg(202) <= s2c(p(201));
	output_reg(201) <= s2c(p(200));
	output_reg(200) <= s2c(p(199));
	output_reg(199) <= s2c(p(198));
	output_reg(198) <= s2c(p(197));
	output_reg(197) <= s2c(p(196));
	output_reg(196) <= s2c(p(195));
	output_reg(195) <= s2c(p(194));
	output_reg(194) <= s2c(p(193));
	output_reg(193) <= s2c(p(192));
	output_reg(192) <= s2c(p(191));
	output_reg(191) <= s2c(p(190));
	output_reg(190) <= s2c(p(189));
	output_reg(189) <= s2c(p(188));
	output_reg(188) <= s2c(p(187));
	output_reg(187) <= s2c(p(186));
	output_reg(186) <= s2c(p(185));
	output_reg(185) <= s2c(p(184));
	output_reg(184) <= s2c(p(183));
	output_reg(183) <= s2c(p(182));
	output_reg(182) <= s2c(p(181));
	output_reg(181) <= s2c(p(180));
	output_reg(180) <= s2c(p(179));
	output_reg(179) <= s2c(p(178));
	output_reg(178) <= s2c(p(177));
	output_reg(177) <= s2c(p(176));
	output_reg(176) <= s2c(p(175));
	output_reg(175) <= s2c(p(174));
	output_reg(174) <= s2c(p(173));
	output_reg(173) <= s2c(p(172));
	output_reg(172) <= s2c(p(171));
	output_reg(171) <= s2c(p(170));
	output_reg(170) <= s2c(p(169));
	output_reg(169) <= s2c(p(168));
	output_reg(168) <= s2c(p(167));
	output_reg(167) <= s2c(p(166));
	output_reg(166) <= s2c(p(165));
	output_reg(165) <= s2c(p(164));
	output_reg(164) <= s2c(p(163));
	output_reg(163) <= s2c(p(162));
	output_reg(162) <= s2c(p(161));
	output_reg(161) <= s2c(p(160));
	output_reg(160) <= s2c(p(159));
	output_reg(159) <= s2c(p(158));
	output_reg(158) <= s2c(p(157));
	output_reg(157) <= s2c(p(156));
	output_reg(156) <= s2c(p(155));
	output_reg(155) <= s2c(p(154));
	output_reg(154) <= s2c(p(153));
	output_reg(153) <= s2c(p(152));
	output_reg(152) <= s2c(p(151));
	output_reg(151) <= s2c(p(150));
	output_reg(150) <= s2c(p(149));
	output_reg(149) <= s2c(p(148));
	output_reg(148) <= s2c(p(147));
	output_reg(147) <= s2c(p(146));
	output_reg(146) <= s2c(p(145));
	output_reg(145) <= s2c(p(144));
	output_reg(144) <= s2c(p(143));
	output_reg(143) <= s2c(p(142));
	output_reg(142) <= s2c(p(141));
	output_reg(141) <= s2c(p(140));
	output_reg(140) <= s2c(p(139));
	output_reg(139) <= s2c(p(138));
	output_reg(138) <= s2c(p(137));
	output_reg(137) <= s2c(p(136));
	output_reg(136) <= s2c(p(135));
	output_reg(135) <= s2c(p(134));
	output_reg(134) <= s2c(p(133));
	output_reg(133) <= s2c(p(132));
	output_reg(132) <= s2c(p(131));
	output_reg(131) <= s2c(p(130));
	output_reg(130) <= s2c(p(129));
	output_reg(129) <= s2c(p(128));
	output_reg(128) <= s2c(p(127));
	output_reg(127) <= s2c(p(126));
	output_reg(126) <= s2c(p(125));
	output_reg(125) <= s2c(p(124));
	output_reg(124) <= s2c(p(123));
	output_reg(123) <= s2c(p(122));
	output_reg(122) <= s2c(p(121));
	output_reg(121) <= s2c(p(120));
	output_reg(120) <= s2c(p(119));
	output_reg(119) <= s2c(p(118));
	output_reg(118) <= s2c(p(117));
	output_reg(117) <= s2c(p(116));
	output_reg(116) <= s2c(p(115));
	output_reg(115) <= s2c(p(114));
	output_reg(114) <= s2c(p(113));
	output_reg(113) <= s2c(p(112));
	output_reg(112) <= s2c(p(111));
	output_reg(111) <= s2c(p(110));
	output_reg(110) <= s2c(p(109));
	output_reg(109) <= s2c(p(108));
	output_reg(108) <= s2c(p(107));
	output_reg(107) <= s2c(p(106));
	output_reg(106) <= s2c(p(105));
	output_reg(105) <= s2c(p(104));
	output_reg(104) <= s2c(p(103));
	output_reg(103) <= s2c(p(102));
	output_reg(102) <= s2c(p(101));
	output_reg(101) <= s2c(p(100));
	output_reg(100) <= s2c(p(99));
	output_reg(99) <= s2c(p(98));
	output_reg(98) <= s2c(p(97));
	output_reg(97) <= s2c(p(96));
	output_reg(96) <= s2c(p(95));
	output_reg(95) <= s2c(p(94));
	output_reg(94) <= s2c(p(93));
	output_reg(93) <= s2c(p(92));
	output_reg(92) <= s2c(p(91));
	output_reg(91) <= s2c(p(90));
	output_reg(90) <= s2c(p(89));
	output_reg(89) <= s2c(p(88));
	output_reg(88) <= s2c(p(87));
	output_reg(87) <= s2c(p(86));
	output_reg(86) <= s2c(p(85));
	output_reg(85) <= s2c(p(84));
	output_reg(84) <= s2c(p(83));
	output_reg(83) <= s2c(p(82));
	output_reg(82) <= s2c(p(81));
	output_reg(81) <= s2c(p(80));
	output_reg(80) <= s2c(p(79));
	output_reg(79) <= s2c(p(78));
	output_reg(78) <= s2c(p(77));
	output_reg(77) <= s2c(p(76));
	output_reg(76) <= s2c(p(75));
	output_reg(75) <= s2c(p(74));
	output_reg(74) <= s2c(p(73));
	output_reg(73) <= s2c(p(72));
	output_reg(72) <= s2c(p(71));
	output_reg(71) <= s2c(p(70));
	output_reg(70) <= s2c(p(69));
	output_reg(69) <= s2c(p(68));
	output_reg(68) <= s2c(p(67));
	output_reg(67) <= s2c(p(66));
	output_reg(66) <= s2c(p(65));
	output_reg(65) <= s2c(p(64));
	output_reg(64) <= s2c(p(63));
	output_reg(63) <= s2c(p(62));
	output_reg(62) <= s2c(p(61));
	output_reg(61) <= s2c(p(60));
	output_reg(60) <= s2c(p(59));
	output_reg(59) <= s2c(p(58));
	output_reg(58) <= s2c(p(57));
	output_reg(57) <= s2c(p(56));
	output_reg(56) <= s2c(p(55));
	output_reg(55) <= s2c(p(54));
	output_reg(54) <= s2c(p(53));
	output_reg(53) <= s2c(p(52));
	output_reg(52) <= s2c(p(51));
	output_reg(51) <= s2c(p(50));
	output_reg(50) <= s2c(p(49));
	output_reg(49) <= s2c(p(48));
	output_reg(48) <= s2c(p(47));
	output_reg(47) <= s2c(p(46));
	output_reg(46) <= s2c(p(45));
	output_reg(45) <= s2c(p(44));
	output_reg(44) <= s2c(p(43));
	output_reg(43) <= s2c(p(42));
	output_reg(42) <= s2c(p(41));
	output_reg(41) <= s2c(p(40));
	output_reg(40) <= s2c(p(39));
	output_reg(39) <= s2c(p(38));
	output_reg(38) <= s2c(p(37));
	output_reg(37) <= s2c(p(36));
	output_reg(36) <= s2c(p(35));
	output_reg(35) <= s2c(p(34));
	output_reg(34) <= s2c(p(33));
	output_reg(33) <= s2c(p(32));
	output_reg(32) <= s2c(p(31));
	output_reg(31) <= s2c(p(30));
	output_reg(30) <= s2c(p(29));
	output_reg(29) <= s2c(p(28));
	output_reg(28) <= s2c(p(27));
	output_reg(27) <= s2c(p(26));
	output_reg(26) <= s2c(p(25));
	output_reg(25) <= s2c(p(24));
	output_reg(24) <= s2c(p(23));
	output_reg(23) <= s2c(p(22));
	output_reg(22) <= s2c(p(21));
	output_reg(21) <= s2c(p(20));
	output_reg(20) <= s2c(p(19));
	output_reg(19) <= s2c(p(18));
	output_reg(18) <= s2c(p(17));
	output_reg(17) <= s2c(p(16));
	output_reg(16) <= s2c(p(15));
	output_reg(15) <= s2c(p(14));
	output_reg(14) <= s2c(p(13));
	output_reg(13) <= s2c(p(12));
	output_reg(12) <= s2c(p(11));
	output_reg(11) <= s2c(p(10));
	output_reg(10) <= s2c(p(9));
	output_reg(9) <= s2c(p(8));
	output_reg(8) <= s2c(p(7));
	output_reg(7) <= s2c(p(6));
	output_reg(6) <= s2c(p(5));
	output_reg(5) <= s2c(p(4));
	output_reg(4) <= s2c(p(3));
	output_reg(3) <= s2c(p(2));
	output_reg(2) <= s2c(p(1));
	output_reg(1) <= s2c(p(0));
	output_reg(0) <= s2c(done);
	---------------------------------------------	
END behavioral;